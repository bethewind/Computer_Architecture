module control(s1, s2, sign, sa, addsub, sr);
input s1, s2, sign, sa;
output addsub, sr;

endmodule