module Multiplier_32(a,b,clk,s);

input [31:0]a,b;
input clk;
output [63:0]s;
wire [:0]w;


//stage1
FA F00(a[1],b[0],a[0],b[1],0,b[2],w[0]);
FA F01(a[2],b[0],a[1],b[1],a[0],b[2],w[1]);
FA F02(a[3],b[0],a[2],b[1],a[1],b[2],w[2]);
FA F03(a[4],b[0],a[3],b[1],a[2],b[2],w[3]);
FA F04(a[5],b[0],a[4],b[1],a[3],b[2],w[4]);
FA F05(a[6],b[0],a[5],b[1],a[4],b[2],w[5]);
FA F06(a[7],b[0],a[6],b[1],a[5],b[2],w[6]);
FA F07(a[8],b[0],a[7],b[1],a[6],b[2],w[7]);
FA F08(a[9],b[0],a[8],b[1],a[7],b[2],w[8]);
FA F09(a[10],b[0],a[9],b[1],a[8],b[2],w[9]);
FA F10(a[11],b[0],a[10],b[1],a[9],b[2],w[10]);
FA F11(a[12],b[0],a[11],b[1],a[10],b[2],w[11]);
FA F12(a[13],b[0],a[12],b[1],a[11],b[2],w[12]);
FA F13(a[14],b[0],a[13],b[1],a[12],b[2],w[13]);
FA F14(a[15],b[0],a[14],b[1],a[13],b[2],w[14]);
FA F15(a[16],b[0],a[15],b[1],a[14],b[2],w[15]);
FA F16(a[17],b[0],a[16],b[1],a[15],b[2],w[16]);
FA F17(a[18],b[0],a[17],b[1],a[16],b[2],w[17]);
FA F18(a[19],b[0],a[18],b[1],a[17],b[2],w[18]);
FA F19(a[20],b[0],a[19],b[1],a[18],b[2],w[19]);
FA F20(a[21],b[0],a[20],b[1],a[19],b[2],w[20]);
FA F21(a[22],b[0],a[21],b[1],a[20],b[2],w[21]);
FA F22(a[23],b[0],a[22],b[1],a[21],b[2],w[22]);
FA F23(a[24],b[0],a[23],b[1],a[22],b[2],w[23]);
FA F24(a[25],b[0],a[24],b[1],a[23],b[2],w[24]);
FA F25(a[26],b[0],a[25],b[1],a[24],b[2],w[25]);
FA F26(a[27],b[0],a[26],b[1],a[25],b[2],w[26]);
FA F27(a[28],b[0],a[27],b[1],a[26],b[2],w[27]);
FA F28(a[29],b[0],a[28],b[1],a[27],b[2],w[28]);
FA F29(a[30],b[0],a[29],b[1],a[28],b[2],w[29]);
FA F30(a[31],b[0],a[30],b[1],a[29],b[2],w[30]);
FA F31(0,b[0],a[31],b[1],a[30],b[2],w[31]);

//STAGE2

FA F1(w[],w[],a[],b[],)

endmodule