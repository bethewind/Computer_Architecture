module rightshifter32(M1, shift, out);
input [31:0]M1;
input [4:0]shift;
output [31:0]out;
wire[160:0]w;

//16bit shift
mux m0(M1[0], M1[16], shift[4], w[0]);
mux m1(M1[1], M1[17], shift[4], w[1]);
mux m2(M1[2], M1[18], shift[4], w[2]);
mux m3(M1[3], M1[19], shift[4], w[3]);
mux m4(M1[4], M1[20], shift[4], w[4]);
mux m5(M1[5], M1[21], shift[4], w[5]);
mux m6(M1[6], M1[22], shift[4], w[6]);
mux m7(M1[7], M1[23], shift[4], w[7]);
mux m8(M1[8], M1[24], shift[4], w[8]);
mux m9(M1[9], M1[25], shift[4], w[9]);
mux M10(M1[10], M1[26], shift[4], w[10]);
mux M11(M1[11], M1[27], shift[4], w[11]);
mux M12(M1[12], M1[28], shift[4], w[12]);
mux M13(M1[13], M1[29], shift[4], w[13]);
mux M14(M1[14], M1[30], shift[4], w[14]);
mux M15(M1[15], M1[31], shift[4], w[15]);
mux M16(M1[16], 1'b0, shift[4], w[16]);
mux M17(M1[17], 1'b0, shift[4], w[17]);
mux M18(M1[18], 1'b0, shift[4], w[18]);
mux M19(M1[19], 1'b0, shift[4], w[19]);
mux m20(M1[20], 1'b0, shift[4], w[20]);
mux m21(M1[21], 1'b0, shift[4], w[21]);
mux m22(M1[22], 1'b0, shift[4], w[22]);
mux m23(M1[23], 1'b0, shift[4], w[23]);
mux m24(M1[24], 1'b0, shift[4], w[24]);
mux m25(M1[25], 1'b0, shift[4], w[25]);
mux m26(M1[26], 1'b0, shift[4], w[26]);
mux m27(M1[27], 1'b0, shift[4], w[27]);
mux m28(M1[28], 1'b0, shift[4], w[28]);
mux m29(M1[29], 1'b0, shift[4], w[29]);
mux m30(M1[30], 1'b0, shift[4], w[30]);
mux m31(M1[31], 1'b0, shift[4], w[31]);

//8bit shift
mux m32(w[0], w[8], shift[3], w[32]);
mux m33(w[1], w[9], shift[3], w[33]);
mux m34(w[2], w[10], shift[3], w[34]);
mux m35(w[3], w[11], shift[3], w[35]);
mux m36(w[4], w[12], shift[3], w[36]);
mux m37(w[5], w[13], shift[3], w[37]);
mux m38(w[6], w[14], shift[3], w[38]);
mux m39(w[7], w[15], shift[3], w[39]);
mux m40(w[8], w[16], shift[3], w[40]);
mux m41(w[9], w[17], shift[3], w[41]);
mux m42(w[10], w[18], shift[3], w[42]);
mux m43(w[11], w[19], shift[3], w[43]);
mux m44(w[12], w[20], shift[3], w[44]);
mux m45(w[13], w[21], shift[3], w[45]);
mux m46(w[14], w[22], shift[3], w[46]);
mux m47(w[15], w[23], shift[3], w[47]);
mux m48(w[16], w[24], shift[3], w[48]);
mux m49(w[17], w[25], shift[3], w[49]);
mux m50(w[18], w[26], shift[3], w[50]);
mux m51(w[19], w[27], shift[3], w[51]);
mux m52(w[20], w[28], shift[3], w[52]);
mux m53(w[21], w[29], shift[3], w[53]);
mux m54(w[22], w[30], shift[3], w[54]);
mux m55(w[23], w[31], shift[3], w[55]);
mux m56(w[24], 1'b0, shift[3], w[56]);
mux m57(w[25], 1'b0, shift[3], w[57]);
mux m58(w[26], 1'b0, shift[3], w[58]);
mux m59(w[27], 1'b0, shift[3], w[59]);
mux m60(w[28], 1'b0, shift[3], w[60]);
mux m61(w[29], 1'b0, shift[3], w[61]);
mux m62(w[30], 1'b0, shift[3], w[62]);
mux m63(w[31], 1'b0, shift[3], w[63]);

//4bit shift
mux m64(w[32], w[36], shift[2], w[64]);
mux m65(w[33], w[37], shift[2], w[65]);
mux m66(w[34], w[38], shift[2], w[66]);
mux m67(w[35], w[39], shift[2], w[67]);
mux m68(w[36], w[40], shift[2], w[68]);
mux m69(w[37], w[41], shift[2], w[69]);
mux m70(w[38], w[42], shift[2], w[70]);
mux m71(w[39], w[43], shift[2], w[71]);
mux m72(w[40], w[44], shift[2], w[72]);
mux m73(w[41], w[45], shift[2], w[73]);
mux m74(w[42], w[46], shift[2], w[74]);
mux m75(w[43], w[47], shift[2], w[75]);
mux m76(w[44], w[48], shift[2], w[76]);
mux m77(w[45], w[49], shift[2], w[77]);
mux m78(w[46], w[50], shift[2], w[78]);
mux m79(w[47], w[51], shift[2], w[79]);
mux m80(w[48], w[52], shift[2], w[80]);
mux m81(w[49], w[53], shift[2], w[81]);
mux m82(w[50], w[54], shift[2], w[82]);
mux m83(w[51], w[55], shift[2], w[83]);
mux m84(w[52], w[56], shift[2], w[84]);
mux m85(w[53], w[57], shift[2], w[85]);
mux m86(w[54], w[58], shift[2], w[86]);
mux m87(w[55], w[59], shift[2], w[87]);
mux m88(w[56], w[60], shift[2], w[88]);
mux m89(w[57], w[61], shift[2], w[89]);
mux m90(w[58], w[62], shift[2], w[90]);
mux m91(w[59], w[63], shift[2], w[91]);
mux m92(w[60], 1'b0, shift[2], w[92]);
mux m93(w[61], 1'b0, shift[2], w[93]);
mux m94(w[62], 1'b0, shift[2], w[94]);
mux m95(w[63], 1'b0, shift[2], w[95]);

assign w[127:96] = w[95:64];

//2bit 
mux M128(w[96], w[98], shift[1], w[128]);
mux M129(w[97], w[99], shift[1], w[129]);
mux M130(w[98], w[100], shift[1], w[130]);
mux M131(w[99], w[101], shift[1], w[131]);
mux M132(w[100], w[102], shift[1], w[132]);
mux M133(w[101], w[103], shift[1], w[133]);
mux M134(w[102], w[104], shift[1], w[134]);
mux M135(w[103], w[105], shift[1], w[135]);
mux M136(w[104], w[106], shift[1], w[136]);
mux M137(w[105], w[107], shift[1], w[137]);
mux M138(w[106], w[108], shift[1], w[138]);
mux M139(w[107], w[109], shift[1], w[139]);
mux M140(w[108], w[110], shift[1], w[140]);
mux M141(w[109], w[111], shift[1], w[141]);
mux M142(w[110], w[112], shift[1], w[142]);
mux M143(w[111], w[113], shift[1], w[143]);
mux M144(w[112], w[114], shift[1], w[144]);
mux M145(w[113], w[115], shift[1], w[145]);
mux M146(w[114], w[116], shift[1], w[146]);
mux M147(w[115], w[117], shift[1], w[147]);
mux M148(w[116], w[118], shift[1], w[148]);
mux M149(w[117], w[119], shift[1], w[149]);
mux M150(w[118], w[120], shift[1], w[150]);
mux M151(w[119], w[121], shift[1], w[151]);
mux M152(w[120], w[122], shift[1], w[152]);
mux M153(w[121], w[123], shift[1], w[153]);
mux M154(w[122], w[124], shift[1], w[154]);
mux M155(w[123], w[125], shift[1], w[155]);
mux M156(w[124], w[126], shift[1], w[156]);
mux M157(w[125], w[127], shift[1], w[157]);
mux M158(w[126], 1'b0, shift[1], w[158]);
mux M159(w[127], 1'b0, shift[1], w[159]);


//1bit
mux M160(w[128], w[129], shift[0], out[0]);
mux M161(w[129], w[130], shift[0], out[1]);
mux M162(w[130], w[131], shift[0], out[2]);
mux M163(w[131], w[132], shift[0], out[3]);
mux M164(w[132], w[133], shift[0], out[4]);
mux M165(w[133], w[134], shift[0], out[5]);
mux M166(w[134], w[135], shift[0], out[6]);
mux M167(w[135], w[136], shift[0], out[7]);
mux M168(w[136], w[137], shift[0], out[8]);
mux M169(w[137], w[138], shift[0], out[9]);
mux M170(w[138], w[139], shift[0], out[10]);
mux M171(w[139], w[140], shift[0], out[11]);
mux M172(w[140], w[141], shift[0], out[12]);
mux M173(w[141], w[142], shift[0], out[13]);
mux M174(w[142], w[143], shift[0], out[14]);
mux M175(w[143], w[144], shift[0], out[15]);
mux M176(w[144], w[145], shift[0], out[16]);
mux M177(w[145], w[146], shift[0], out[17]);
mux M178(w[146], w[147], shift[0], out[18]);
mux M179(w[147], w[148], shift[0], out[19]);
mux M180(w[148], w[149], shift[0], out[20]);
mux M181(w[149], w[150], shift[0], out[21]);
mux M182(w[150], w[151], shift[0], out[22]);
mux M183(w[151], w[152], shift[0], out[23]);
mux M184(w[152], w[153], shift[0], out[24]);
mux M185(w[153], w[154], shift[0], out[25]);
mux M186(w[154], w[155], shift[0], out[26]);
mux M187(w[155], w[156], shift[0], out[27]);
mux M188(w[156], w[157], shift[0], out[28]);
mux M189(w[157], w[158], shift[0], out[29]);
mux M190(w[158], w[159], shift[0], out[30]);
mux M191(w[159], 1'b0, shift[0], out[31]);

endmodule