module Cache(x,y,word,counter);
input [11:0]x;
output reg y;
output [7:0]word;
output [2:0]counter;

reg [63:0]cache[63:0];
reg [63:0]MM[511:0];
reg [8:0]tag[63:0];
reg [63:0]buff;
reg flag;
reg [2:0]index;
reg [2:0]pointer;

wire [8:0]t;
wire [2:0]bo;
wire [7:0]temp;

assign t = x[11:3];
assign bo = x[2:0];

initial 
begin

pointer = 3'b000;

flag = 0;
index = 3'b000;


cache[0] = 64'd0;
cache[1] = 64'd0;
cache[2] = 64'd0;
cache[3] = 64'd0;
cache[4] = 64'd0;
cache[5] = 64'd0;
cache[6] = 64'd0;
cache[7] = 64'd0;


tag[0] = 9'd0;
tag[1] = 9'd0;
tag[2] = 9'd0;
tag[3] = 9'd0;
tag[4] = 9'd16;
tag[5] = 9'd0;
tag[6] = 9'd0;
tag[7] = 9'd0;


MM[0] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
MM[1] = 64'b1111111111111111111111111111111111111111111111111111111111111110;
MM[2] = 64'b1111111111111111111111111111111111111111111111111111111111111101;
MM[3] = 64'b1111111111111111111111111111111111111111111111111111111111111100;
MM[4] = 64'b1111111111111111111111111111111111111111111111111111111111111011;
MM[5] = 64'b1111111111111111111111111111111111111111111111111111111111111010;
MM[6] = 64'b1111111111111111111111111111111111111111111111111111111111111001;
MM[7] = 64'b1111111111111111111111111111111111111111111111111111111111111000;
MM[8] = 64'b1111111111111111111111111111111111111111111111111111111111110111;
MM[9] = 64'b1111111111111111111111111111111111111111111111111111111111110110;
MM[10] = 64'b1111111111111111111111111111111111111111111111111111111111110101;
MM[11] = 64'b1111111111111111111111111111111111111111111111111111111111110100;
MM[12] = 64'b1111111111111111111111111111111111111111111111111111111111110011;
MM[13] = 64'b1111111111111111111111111111111111111111111111111111111111110010;
MM[14] = 64'b1111111111111111111111111111111111111111111111111111111111110001;
MM[15] = 64'b1111111111111111111111111111111111111111111111111111111111110000;
MM[16] = 64'b1111111111111111111111111111111111111111111111111111111111101111;
MM[17] = 64'b1111111111111111111111111111111111111111111111111111111111101110;
MM[18] = 64'b1111111111111111111111111111111111111111111111111111111111101101;
MM[19] = 64'b1111111111111111111111111111111111111111111111111111111111101100;
MM[20] = 64'b1111111111111111111111111111111111111111111111111111111111101011;
MM[21] = 64'b1111111111111111111111111111111111111111111111111111111111101010;
MM[22] = 64'b1111111111111111111111111111111111111111111111111111111111101001;
MM[23] = 64'b1111111111111111111111111111111111111111111111111111111111101000;
MM[24] = 64'b1111111111111111111111111111111111111111111111111111111111100111;
MM[25] = 64'b1111111111111111111111111111111111111111111111111111111111100110;
MM[26] = 64'b1111111111111111111111111111111111111111111111111111111111100101;
MM[27] = 64'b1111111111111111111111111111111111111111111111111111111111100100;
MM[28] = 64'b1111111111111111111111111111111111111111111111111111111111100011;
MM[29] = 64'b1111111111111111111111111111111111111111111111111111111111100010;
MM[30] = 64'b1111111111111111111111111111111111111111111111111111111111100001;
MM[31] = 64'b1111111111111111111111111111111111111111111111111111111111100000;
MM[32] = 64'b1111111111111111111111111111111111111111111111111111111111011111;
MM[33] = 64'b1111111111111111111111111111111111111111111111111111111111011110;
MM[34] = 64'b1111111111111111111111111111111111111111111111111111111111011101;
MM[35] = 64'b1111111111111111111111111111111111111111111111111111111111011100;
MM[36] = 64'b1111111111111111111111111111111111111111111111111111111111011011;
MM[37] = 64'b1111111111111111111111111111111111111111111111111111111111011010;
MM[38] = 64'b1111111111111111111111111111111111111111111111111111111111011001;
MM[39] = 64'b1111111111111111111111111111111111111111111111111111111111011000;
MM[40] = 64'b1111111111111111111111111111111111111111111111111111111111010111;
MM[41] = 64'b1111111111111111111111111111111111111111111111111111111111010110;
MM[42] = 64'b1111111111111111111111111111111111111111111111111111111111010101;
MM[43] = 64'b1111111111111111111111111111111111111111111111111111111111010100;
MM[44] = 64'b1111111111111111111111111111111111111111111111111111111111010011;
MM[45] = 64'b1111111111111111111111111111111111111111111111111111111111010010;
MM[46] = 64'b1111111111111111111111111111111111111111111111111111111111010001;
MM[47] = 64'b1111111111111111111111111111111111111111111111111111111111010000;
MM[48] = 64'b1111111111111111111111111111111111111111111111111111111111001111;
MM[49] = 64'b1111111111111111111111111111111111111111111111111111111111001110;
MM[50] = 64'b1111111111111111111111111111111111111111111111111111111111001101;
MM[51] = 64'b1111111111111111111111111111111111111111111111111111111111001100;
MM[52] = 64'b1111111111111111111111111111111111111111111111111111111111001011;
MM[53] = 64'b1111111111111111111111111111111111111111111111111111111111001010;
MM[54] = 64'b1111111111111111111111111111111111111111111111111111111111001001;
MM[55] = 64'b1111111111111111111111111111111111111111111111111111111111001000;
MM[56] = 64'b1111111111111111111111111111111111111111111111111111111111000111;
MM[57] = 64'b1111111111111111111111111111111111111111111111111111111111000110;
MM[58] = 64'b1111111111111111111111111111111111111111111111111111111111000101;
MM[59] = 64'b1111111111111111111111111111111111111111111111111111111111000100;
MM[60] = 64'b1111111111111111111111111111111111111111111111111111111111000011;
MM[61] = 64'b1111111111111111111111111111111111111111111111111111111111000010;
MM[62] = 64'b1111111111111111111111111111111111111111111111111111111111000001;
MM[63] = 64'b1111111111111111111111111111111111111111111111111111111111000000;
MM[64] = 64'b1111111111111111111111111111111111111111111111111111111110111111;
MM[65] = 64'b1111111111111111111111111111111111111111111111111111111110111110;
MM[66] = 64'b1111111111111111111111111111111111111111111111111111111110111101;
MM[67] = 64'b1111111111111111111111111111111111111111111111111111111110111100;
MM[68] = 64'b1111111111111111111111111111111111111111111111111111111110111011;
MM[69] = 64'b1111111111111111111111111111111111111111111111111111111110111010;
MM[70] = 64'b1111111111111111111111111111111111111111111111111111111110111001;
MM[71] = 64'b1111111111111111111111111111111111111111111111111111111110111000;
MM[72] = 64'b1111111111111111111111111111111111111111111111111111111110110111;
MM[73] = 64'b1111111111111111111111111111111111111111111111111111111110110110;
MM[74] = 64'b1111111111111111111111111111111111111111111111111111111110110101;
MM[75] = 64'b1111111111111111111111111111111111111111111111111111111110110100;
MM[76] = 64'b1111111111111111111111111111111111111111111111111111111110110011;
MM[77] = 64'b1111111111111111111111111111111111111111111111111111111110110010;
MM[78] = 64'b1111111111111111111111111111111111111111111111111111111110110001;
MM[79] = 64'b1111111111111111111111111111111111111111111111111111111110110000;
MM[80] = 64'b1111111111111111111111111111111111111111111111111111111110101111;
MM[81] = 64'b1111111111111111111111111111111111111111111111111111111110101110;
MM[82] = 64'b1111111111111111111111111111111111111111111111111111111110101101;
MM[83] = 64'b1111111111111111111111111111111111111111111111111111111110101100;
MM[84] = 64'b1111111111111111111111111111111111111111111111111111111110101011;
MM[85] = 64'b1111111111111111111111111111111111111111111111111111111110101010;
MM[86] = 64'b1111111111111111111111111111111111111111111111111111111110101001;
MM[87] = 64'b1111111111111111111111111111111111111111111111111111111110101000;
MM[88] = 64'b1111111111111111111111111111111111111111111111111111111110100111;
MM[89] = 64'b1111111111111111111111111111111111111111111111111111111110100110;
MM[90] = 64'b1111111111111111111111111111111111111111111111111111111110100101;
MM[91] = 64'b1111111111111111111111111111111111111111111111111111111110100100;
MM[92] = 64'b1111111111111111111111111111111111111111111111111111111110100011;
MM[93] = 64'b1111111111111111111111111111111111111111111111111111111110100010;
MM[94] = 64'b1111111111111111111111111111111111111111111111111111111110100001;
MM[95] = 64'b1111111111111111111111111111111111111111111111111111111110100000;
MM[96] = 64'b1111111111111111111111111111111111111111111111111111111110011111;
MM[97] = 64'b1111111111111111111111111111111111111111111111111111111110011110;
MM[98] = 64'b1111111111111111111111111111111111111111111111111111111110011101;
MM[99] = 64'b1111111111111111111111111111111111111111111111111111111110011100;
MM[100] = 64'b1111111111111111111111111111111111111111111111111111111110011011;
MM[101] = 64'b1111111111111111111111111111111111111111111111111111111110011010;
MM[102] = 64'b1111111111111111111111111111111111111111111111111111111110011001;
MM[103] = 64'b1111111111111111111111111111111111111111111111111111111110011000;
MM[104] = 64'b1111111111111111111111111111111111111111111111111111111110010111;
MM[105] = 64'b1111111111111111111111111111111111111111111111111111111110010110;
MM[106] = 64'b1111111111111111111111111111111111111111111111111111111110010101;
MM[107] = 64'b1111111111111111111111111111111111111111111111111111111110010100;
MM[108] = 64'b1111111111111111111111111111111111111111111111111111111110010011;
MM[109] = 64'b1111111111111111111111111111111111111111111111111111111110010010;
MM[110] = 64'b1111111111111111111111111111111111111111111111111111111110010001;
MM[111] = 64'b1111111111111111111111111111111111111111111111111111111110010000;
MM[112] = 64'b1111111111111111111111111111111111111111111111111111111110001111;
MM[113] = 64'b1111111111111111111111111111111111111111111111111111111110001110;
MM[114] = 64'b1111111111111111111111111111111111111111111111111111111110001101;
MM[115] = 64'b1111111111111111111111111111111111111111111111111111111110001100;
MM[116] = 64'b1111111111111111111111111111111111111111111111111111111110001011;
MM[117] = 64'b1111111111111111111111111111111111111111111111111111111110001010;
MM[118] = 64'b1111111111111111111111111111111111111111111111111111111110001001;
MM[119] = 64'b1111111111111111111111111111111111111111111111111111111110001000;
MM[120] = 64'b1111111111111111111111111111111111111111111111111111111110000111;
MM[121] = 64'b1111111111111111111111111111111111111111111111111111111110000110;
MM[122] = 64'b1111111111111111111111111111111111111111111111111111111110000101;
MM[123] = 64'b1111111111111111111111111111111111111111111111111111111110000100;
MM[124] = 64'b1111111111111111111111111111111111111111111111111111111110000011;
MM[125] = 64'b1111111111111111111111111111111111111111111111111111111110000010;
MM[126] = 64'b1111111111111111111111111111111111111111111111111111111110000001;
MM[127] = 64'b1111111111111111111111111111111111111111111111111111111110000000;
MM[128] = 64'b1111111111111111111111111111111111111111111111111111111101111111;
MM[129] = 64'b1111111111111111111111111111111111111111111111111111111101111110;
MM[130] = 64'b1111111111111111111111111111111111111111111111111111111101111101;
MM[131] = 64'b1111111111111111111111111111111111111111111111111111111101111100;
MM[132] = 64'b1111111111111111111111111111111111111111111111111111111101111011;
MM[133] = 64'b1111111111111111111111111111111111111111111111111111111101111010;
MM[134] = 64'b1111111111111111111111111111111111111111111111111111111101111001;
MM[135] = 64'b1111111111111111111111111111111111111111111111111111111101111000;
MM[136] = 64'b1111111111111111111111111111111111111111111111111111111101110111;
MM[137] = 64'b1111111111111111111111111111111111111111111111111111111101110110;
MM[138] = 64'b1111111111111111111111111111111111111111111111111111111101110101;
MM[139] = 64'b1111111111111111111111111111111111111111111111111111111101110100;
MM[140] = 64'b1111111111111111111111111111111111111111111111111111111101110011;
MM[141] = 64'b1111111111111111111111111111111111111111111111111111111101110010;
MM[142] = 64'b1111111111111111111111111111111111111111111111111111111101110001;
MM[143] = 64'b1111111111111111111111111111111111111111111111111111111101110000;
MM[144] = 64'b1111111111111111111111111111111111111111111111111111111101101111;
MM[145] = 64'b1111111111111111111111111111111111111111111111111111111101101110;
MM[146] = 64'b1111111111111111111111111111111111111111111111111111111101101101;
MM[147] = 64'b1111111111111111111111111111111111111111111111111111111101101100;
MM[148] = 64'b1111111111111111111111111111111111111111111111111111111101101011;
MM[149] = 64'b1111111111111111111111111111111111111111111111111111111101101010;
MM[150] = 64'b1111111111111111111111111111111111111111111111111111111101101001;
MM[151] = 64'b1111111111111111111111111111111111111111111111111111111101101000;
MM[152] = 64'b1111111111111111111111111111111111111111111111111111111101100111;
MM[153] = 64'b1111111111111111111111111111111111111111111111111111111101100110;
MM[154] = 64'b1111111111111111111111111111111111111111111111111111111101100101;
MM[155] = 64'b1111111111111111111111111111111111111111111111111111111101100100;
MM[156] = 64'b1111111111111111111111111111111111111111111111111111111101100011;
MM[157] = 64'b1111111111111111111111111111111111111111111111111111111101100010;
MM[158] = 64'b1111111111111111111111111111111111111111111111111111111101100001;
MM[159] = 64'b1111111111111111111111111111111111111111111111111111111101100000;
MM[160] = 64'b1111111111111111111111111111111111111111111111111111111101011111;
MM[161] = 64'b1111111111111111111111111111111111111111111111111111111101011110;
MM[162] = 64'b1111111111111111111111111111111111111111111111111111111101011101;
MM[163] = 64'b1111111111111111111111111111111111111111111111111111111101011100;
MM[164] = 64'b1111111111111111111111111111111111111111111111111111111101011011;
MM[165] = 64'b1111111111111111111111111111111111111111111111111111111101011010;
MM[166] = 64'b1111111111111111111111111111111111111111111111111111111101011001;
MM[167] = 64'b1111111111111111111111111111111111111111111111111111111101011000;
MM[168] = 64'b1111111111111111111111111111111111111111111111111111111101010111;
MM[169] = 64'b1111111111111111111111111111111111111111111111111111111101010110;
MM[170] = 64'b1111111111111111111111111111111111111111111111111111111101010101;
MM[171] = 64'b1111111111111111111111111111111111111111111111111111111101010100;
MM[172] = 64'b1111111111111111111111111111111111111111111111111111111101010011;
MM[173] = 64'b1111111111111111111111111111111111111111111111111111111101010010;
MM[174] = 64'b1111111111111111111111111111111111111111111111111111111101010001;
MM[175] = 64'b1111111111111111111111111111111111111111111111111111111101010000;
MM[176] = 64'b1111111111111111111111111111111111111111111111111111111101001111;
MM[177] = 64'b1111111111111111111111111111111111111111111111111111111101001110;
MM[178] = 64'b1111111111111111111111111111111111111111111111111111111101001101;
MM[179] = 64'b1111111111111111111111111111111111111111111111111111111101001100;
MM[180] = 64'b1111111111111111111111111111111111111111111111111111111101001011;
MM[181] = 64'b1111111111111111111111111111111111111111111111111111111101001010;
MM[182] = 64'b1111111111111111111111111111111111111111111111111111111101001001;
MM[183] = 64'b1111111111111111111111111111111111111111111111111111111101001000;
MM[184] = 64'b1111111111111111111111111111111111111111111111111111111101000111;
MM[185] = 64'b1111111111111111111111111111111111111111111111111111111101000110;
MM[186] = 64'b1111111111111111111111111111111111111111111111111111111101000101;
MM[187] = 64'b1111111111111111111111111111111111111111111111111111111101000100;
MM[188] = 64'b1111111111111111111111111111111111111111111111111111111101000011;
MM[189] = 64'b1111111111111111111111111111111111111111111111111111111101000010;
MM[190] = 64'b1111111111111111111111111111111111111111111111111111111101000001;
MM[191] = 64'b1111111111111111111111111111111111111111111111111111111101000000;
MM[192] = 64'b1111111111111111111111111111111111111111111111111111111100111111;
MM[193] = 64'b1111111111111111111111111111111111111111111111111111111100111110;
MM[194] = 64'b1111111111111111111111111111111111111111111111111111111100111101;
MM[195] = 64'b1111111111111111111111111111111111111111111111111111111100111100;
MM[196] = 64'b1111111111111111111111111111111111111111111111111111111100111011;
MM[197] = 64'b1111111111111111111111111111111111111111111111111111111100111010;
MM[198] = 64'b1111111111111111111111111111111111111111111111111111111100111001;
MM[199] = 64'b1111111111111111111111111111111111111111111111111111111100111000;
MM[200] = 64'b1111111111111111111111111111111111111111111111111111111100110111;
MM[201] = 64'b1111111111111111111111111111111111111111111111111111111100110110;
MM[202] = 64'b1111111111111111111111111111111111111111111111111111111100110101;
MM[203] = 64'b1111111111111111111111111111111111111111111111111111111100110100;
MM[204] = 64'b1111111111111111111111111111111111111111111111111111111100110011;
MM[205] = 64'b1111111111111111111111111111111111111111111111111111111100110010;
MM[206] = 64'b1111111111111111111111111111111111111111111111111111111100110001;
MM[207] = 64'b1111111111111111111111111111111111111111111111111111111100110000;
MM[208] = 64'b1111111111111111111111111111111111111111111111111111111100101111;
MM[209] = 64'b1111111111111111111111111111111111111111111111111111111100101110;
MM[210] = 64'b1111111111111111111111111111111111111111111111111111111100101101;
MM[211] = 64'b1111111111111111111111111111111111111111111111111111111100101100;
MM[212] = 64'b1111111111111111111111111111111111111111111111111111111100101011;
MM[213] = 64'b1111111111111111111111111111111111111111111111111111111100101010;
MM[214] = 64'b1111111111111111111111111111111111111111111111111111111100101001;
MM[215] = 64'b1111111111111111111111111111111111111111111111111111111100101000;
MM[216] = 64'b1111111111111111111111111111111111111111111111111111111100100111;
MM[217] = 64'b1111111111111111111111111111111111111111111111111111111100100110;
MM[218] = 64'b1111111111111111111111111111111111111111111111111111111100100101;
MM[219] = 64'b1111111111111111111111111111111111111111111111111111111100100100;
MM[220] = 64'b1111111111111111111111111111111111111111111111111111111100100011;
MM[221] = 64'b1111111111111111111111111111111111111111111111111111111100100010;
MM[222] = 64'b1111111111111111111111111111111111111111111111111111111100100001;
MM[223] = 64'b1111111111111111111111111111111111111111111111111111111100100000;
MM[224] = 64'b1111111111111111111111111111111111111111111111111111111100011111;
MM[225] = 64'b1111111111111111111111111111111111111111111111111111111100011110;
MM[226] = 64'b1111111111111111111111111111111111111111111111111111111100011101;
MM[227] = 64'b1111111111111111111111111111111111111111111111111111111100011100;
MM[228] = 64'b1111111111111111111111111111111111111111111111111111111100011011;
MM[229] = 64'b1111111111111111111111111111111111111111111111111111111100011010;
MM[230] = 64'b1111111111111111111111111111111111111111111111111111111100011001;
MM[231] = 64'b1111111111111111111111111111111111111111111111111111111100011000;
MM[232] = 64'b1111111111111111111111111111111111111111111111111111111100010111;
MM[233] = 64'b1111111111111111111111111111111111111111111111111111111100010110;
MM[234] = 64'b1111111111111111111111111111111111111111111111111111111100010101;
MM[235] = 64'b1111111111111111111111111111111111111111111111111111111100010100;
MM[236] = 64'b1111111111111111111111111111111111111111111111111111111100010011;
MM[237] = 64'b1111111111111111111111111111111111111111111111111111111100010010;
MM[238] = 64'b1111111111111111111111111111111111111111111111111111111100010001;
MM[239] = 64'b1111111111111111111111111111111111111111111111111111111100010000;
MM[240] = 64'b1111111111111111111111111111111111111111111111111111111100001111;
MM[241] = 64'b1111111111111111111111111111111111111111111111111111111100001110;
MM[242] = 64'b1111111111111111111111111111111111111111111111111111111100001101;
MM[243] = 64'b1111111111111111111111111111111111111111111111111111111100001100;
MM[244] = 64'b1111111111111111111111111111111111111111111111111111111100001011;
MM[245] = 64'b1111111111111111111111111111111111111111111111111111111100001010;
MM[246] = 64'b1111111111111111111111111111111111111111111111111111111100001001;
MM[247] = 64'b1111111111111111111111111111111111111111111111111111111100001000;
MM[248] = 64'b1111111111111111111111111111111111111111111111111111111100000111;
MM[249] = 64'b1111111111111111111111111111111111111111111111111111111100000110;
MM[250] = 64'b1111111111111111111111111111111111111111111111111111111100000101;
MM[251] = 64'b1111111111111111111111111111111111111111111111111111111100000100;
MM[252] = 64'b1111111111111111111111111111111111111111111111111111111100000011;
MM[253] = 64'b1111111111111111111111111111111111111111111111111111111100000010;
MM[254] = 64'b1111111111111111111111111111111111111111111111111111111100000001;
MM[255] = 64'b1111111111111111111111111111111111111111111111111111111100000000;
MM[256] = 64'b1111111111111111111111111111111111111111111111111111111011111111;
MM[257] = 64'b1111111111111111111111111111111111111111111111111111111011111110;
MM[258] = 64'b1111111111111111111111111111111111111111111111111111111011111101;
MM[259] = 64'b1111111111111111111111111111111111111111111111111111111011111100;
MM[260] = 64'b1111111111111111111111111111111111111111111111111111111011111011;
MM[261] = 64'b1111111111111111111111111111111111111111111111111111111011111010;
MM[262] = 64'b1111111111111111111111111111111111111111111111111111111011111001;
MM[263] = 64'b1111111111111111111111111111111111111111111111111111111011111000;
MM[264] = 64'b1111111111111111111111111111111111111111111111111111111011110111;
MM[265] = 64'b1111111111111111111111111111111111111111111111111111111011110110;
MM[266] = 64'b1111111111111111111111111111111111111111111111111111111011110101;
MM[267] = 64'b1111111111111111111111111111111111111111111111111111111011110100;
MM[268] = 64'b1111111111111111111111111111111111111111111111111111111011110011;
MM[269] = 64'b1111111111111111111111111111111111111111111111111111111011110010;
MM[270] = 64'b1111111111111111111111111111111111111111111111111111111011110001;
MM[271] = 64'b1111111111111111111111111111111111111111111111111111111011110000;
MM[272] = 64'b1111111111111111111111111111111111111111111111111111111011101111;
MM[273] = 64'b1111111111111111111111111111111111111111111111111111111011101110;
MM[274] = 64'b1111111111111111111111111111111111111111111111111111111011101101;
MM[275] = 64'b1111111111111111111111111111111111111111111111111111111011101100;
MM[276] = 64'b1111111111111111111111111111111111111111111111111111111011101011;
MM[277] = 64'b1111111111111111111111111111111111111111111111111111111011101010;
MM[278] = 64'b1111111111111111111111111111111111111111111111111111111011101001;
MM[279] = 64'b1111111111111111111111111111111111111111111111111111111011101000;
MM[280] = 64'b1111111111111111111111111111111111111111111111111111111011100111;
MM[281] = 64'b1111111111111111111111111111111111111111111111111111111011100110;
MM[282] = 64'b1111111111111111111111111111111111111111111111111111111011100101;
MM[283] = 64'b1111111111111111111111111111111111111111111111111111111011100100;
MM[284] = 64'b1111111111111111111111111111111111111111111111111111111011100011;
MM[285] = 64'b1111111111111111111111111111111111111111111111111111111011100010;
MM[286] = 64'b1111111111111111111111111111111111111111111111111111111011100001;
MM[287] = 64'b1111111111111111111111111111111111111111111111111111111011100000;
MM[288] = 64'b1111111111111111111111111111111111111111111111111111111011011111;
MM[289] = 64'b1111111111111111111111111111111111111111111111111111111011011110;
MM[290] = 64'b1111111111111111111111111111111111111111111111111111111011011101;
MM[291] = 64'b1111111111111111111111111111111111111111111111111111111011011100;
MM[292] = 64'b1111111111111111111111111111111111111111111111111111111011011011;
MM[293] = 64'b1111111111111111111111111111111111111111111111111111111011011010;
MM[294] = 64'b1111111111111111111111111111111111111111111111111111111011011001;
MM[295] = 64'b1111111111111111111111111111111111111111111111111111111011011000;
MM[296] = 64'b1111111111111111111111111111111111111111111111111111111011010111;
MM[297] = 64'b1111111111111111111111111111111111111111111111111111111011010110;
MM[298] = 64'b1111111111111111111111111111111111111111111111111111111011010101;
MM[299] = 64'b1111111111111111111111111111111111111111111111111111111011010100;
MM[300] = 64'b1111111111111111111111111111111111111111111111111111111011010011;
MM[301] = 64'b1111111111111111111111111111111111111111111111111111111011010010;
MM[302] = 64'b1111111111111111111111111111111111111111111111111111111011010001;
MM[303] = 64'b1111111111111111111111111111111111111111111111111111111011010000;
MM[304] = 64'b1111111111111111111111111111111111111111111111111111111011001111;
MM[305] = 64'b1111111111111111111111111111111111111111111111111111111011001110;
MM[306] = 64'b1111111111111111111111111111111111111111111111111111111011001101;
MM[307] = 64'b1111111111111111111111111111111111111111111111111111111011001100;
MM[308] = 64'b1111111111111111111111111111111111111111111111111111111011001011;
MM[309] = 64'b1111111111111111111111111111111111111111111111111111111011001010;
MM[310] = 64'b1111111111111111111111111111111111111111111111111111111011001001;
MM[311] = 64'b1111111111111111111111111111111111111111111111111111111011001000;
MM[312] = 64'b1111111111111111111111111111111111111111111111111111111011000111;
MM[313] = 64'b1111111111111111111111111111111111111111111111111111111011000110;
MM[314] = 64'b1111111111111111111111111111111111111111111111111111111011000101;
MM[315] = 64'b1111111111111111111111111111111111111111111111111111111011000100;
MM[316] = 64'b1111111111111111111111111111111111111111111111111111111011000011;
MM[317] = 64'b1111111111111111111111111111111111111111111111111111111011000010;
MM[318] = 64'b1111111111111111111111111111111111111111111111111111111011000001;
MM[319] = 64'b1111111111111111111111111111111111111111111111111111111011000000;
MM[320] = 64'b1111111111111111111111111111111111111111111111111111111010111111;
MM[321] = 64'b1111111111111111111111111111111111111111111111111111111010111110;
MM[322] = 64'b1111111111111111111111111111111111111111111111111111111010111101;
MM[323] = 64'b1111111111111111111111111111111111111111111111111111111010111100;
MM[324] = 64'b1111111111111111111111111111111111111111111111111111111010111011;
MM[325] = 64'b1111111111111111111111111111111111111111111111111111111010111010;
MM[326] = 64'b1111111111111111111111111111111111111111111111111111111010111001;
MM[327] = 64'b1111111111111111111111111111111111111111111111111111111010111000;
MM[328] = 64'b1111111111111111111111111111111111111111111111111111111010110111;
MM[329] = 64'b1111111111111111111111111111111111111111111111111111111010110110;
MM[330] = 64'b1111111111111111111111111111111111111111111111111111111010110101;
MM[331] = 64'b1111111111111111111111111111111111111111111111111111111010110100;
MM[332] = 64'b1111111111111111111111111111111111111111111111111111111010110011;
MM[333] = 64'b1111111111111111111111111111111111111111111111111111111010110010;
MM[334] = 64'b1111111111111111111111111111111111111111111111111111111010110001;
MM[335] = 64'b1111111111111111111111111111111111111111111111111111111010110000;
MM[336] = 64'b1111111111111111111111111111111111111111111111111111111010101111;
MM[337] = 64'b1111111111111111111111111111111111111111111111111111111010101110;
MM[338] = 64'b1111111111111111111111111111111111111111111111111111111010101101;
MM[339] = 64'b1111111111111111111111111111111111111111111111111111111010101100;
MM[340] = 64'b1111111111111111111111111111111111111111111111111111111010101011;
MM[341] = 64'b1111111111111111111111111111111111111111111111111111111010101010;
MM[342] = 64'b1111111111111111111111111111111111111111111111111111111010101001;
MM[343] = 64'b1111111111111111111111111111111111111111111111111111111010101000;
MM[344] = 64'b1111111111111111111111111111111111111111111111111111111010100111;
MM[345] = 64'b1111111111111111111111111111111111111111111111111111111010100110;
MM[346] = 64'b1111111111111111111111111111111111111111111111111111111010100101;
MM[347] = 64'b1111111111111111111111111111111111111111111111111111111010100100;
MM[348] = 64'b1111111111111111111111111111111111111111111111111111111010100011;
MM[349] = 64'b1111111111111111111111111111111111111111111111111111111010100010;
MM[350] = 64'b1111111111111111111111111111111111111111111111111111111010100001;
MM[351] = 64'b1111111111111111111111111111111111111111111111111111111010100000;
MM[352] = 64'b1111111111111111111111111111111111111111111111111111111010011111;
MM[353] = 64'b1111111111111111111111111111111111111111111111111111111010011110;
MM[354] = 64'b1111111111111111111111111111111111111111111111111111111010011101;
MM[355] = 64'b1111111111111111111111111111111111111111111111111111111010011100;
MM[356] = 64'b1111111111111111111111111111111111111111111111111111111010011011;
MM[357] = 64'b1111111111111111111111111111111111111111111111111111111010011010;
MM[358] = 64'b1111111111111111111111111111111111111111111111111111111010011001;
MM[359] = 64'b1111111111111111111111111111111111111111111111111111111010011000;
MM[360] = 64'b1111111111111111111111111111111111111111111111111111111010010111;
MM[361] = 64'b1111111111111111111111111111111111111111111111111111111010010110;
MM[362] = 64'b1111111111111111111111111111111111111111111111111111111010010101;
MM[363] = 64'b1111111111111111111111111111111111111111111111111111111010010100;
MM[364] = 64'b1111111111111111111111111111111111111111111111111111111010010011;
MM[365] = 64'b1111111111111111111111111111111111111111111111111111111010010010;
MM[366] = 64'b1111111111111111111111111111111111111111111111111111111010010001;
MM[367] = 64'b1111111111111111111111111111111111111111111111111111111010010000;
MM[368] = 64'b1111111111111111111111111111111111111111111111111111111010001111;
MM[369] = 64'b1111111111111111111111111111111111111111111111111111111010001110;
MM[370] = 64'b1111111111111111111111111111111111111111111111111111111010001101;
MM[371] = 64'b1111111111111111111111111111111111111111111111111111111010001100;
MM[372] = 64'b1111111111111111111111111111111111111111111111111111111010001011;
MM[373] = 64'b1111111111111111111111111111111111111111111111111111111010001010;
MM[374] = 64'b1111111111111111111111111111111111111111111111111111111010001001;
MM[375] = 64'b1111111111111111111111111111111111111111111111111111111010001000;
MM[376] = 64'b1111111111111111111111111111111111111111111111111111111010000111;
MM[377] = 64'b1111111111111111111111111111111111111111111111111111111010000110;
MM[378] = 64'b1111111111111111111111111111111111111111111111111111111010000101;
MM[379] = 64'b1111111111111111111111111111111111111111111111111111111010000100;
MM[380] = 64'b1111111111111111111111111111111111111111111111111111111010000011;
MM[381] = 64'b1111111111111111111111111111111111111111111111111111111010000010;
MM[382] = 64'b1111111111111111111111111111111111111111111111111111111010000001;
MM[383] = 64'b1111111111111111111111111111111111111111111111111111111010000000;
MM[384] = 64'b1111111111111111111111111111111111111111111111111111111001111111;
MM[385] = 64'b1111111111111111111111111111111111111111111111111111111001111110;
MM[386] = 64'b1111111111111111111111111111111111111111111111111111111001111101;
MM[387] = 64'b1111111111111111111111111111111111111111111111111111111001111100;
MM[388] = 64'b1111111111111111111111111111111111111111111111111111111001111011;
MM[389] = 64'b1111111111111111111111111111111111111111111111111111111001111010;
MM[390] = 64'b1111111111111111111111111111111111111111111111111111111001111001;
MM[391] = 64'b1111111111111111111111111111111111111111111111111111111001111000;
MM[392] = 64'b1111111111111111111111111111111111111111111111111111111001110111;
MM[393] = 64'b1111111111111111111111111111111111111111111111111111111001110110;
MM[394] = 64'b1111111111111111111111111111111111111111111111111111111001110101;
MM[395] = 64'b1111111111111111111111111111111111111111111111111111111001110100;
MM[396] = 64'b1111111111111111111111111111111111111111111111111111111001110011;
MM[397] = 64'b1111111111111111111111111111111111111111111111111111111001110010;
MM[398] = 64'b1111111111111111111111111111111111111111111111111111111001110001;
MM[399] = 64'b1111111111111111111111111111111111111111111111111111111001110000;
MM[400] = 64'b1111111111111111111111111111111111111111111111111111111001101111;
MM[401] = 64'b1111111111111111111111111111111111111111111111111111111001101110;
MM[402] = 64'b1111111111111111111111111111111111111111111111111111111001101101;
MM[403] = 64'b1111111111111111111111111111111111111111111111111111111001101100;
MM[404] = 64'b1111111111111111111111111111111111111111111111111111111001101011;
MM[405] = 64'b1111111111111111111111111111111111111111111111111111111001101010;
MM[406] = 64'b1111111111111111111111111111111111111111111111111111111001101001;
MM[407] = 64'b1111111111111111111111111111111111111111111111111111111001101000;
MM[408] = 64'b1111111111111111111111111111111111111111111111111111111001100111;
MM[409] = 64'b1111111111111111111111111111111111111111111111111111111001100110;
MM[410] = 64'b1111111111111111111111111111111111111111111111111111111001100101;
MM[411] = 64'b1111111111111111111111111111111111111111111111111111111001100100;
MM[412] = 64'b1111111111111111111111111111111111111111111111111111111001100011;
MM[413] = 64'b1111111111111111111111111111111111111111111111111111111001100010;
MM[414] = 64'b1111111111111111111111111111111111111111111111111111111001100001;
MM[415] = 64'b1111111111111111111111111111111111111111111111111111111001100000;
MM[416] = 64'b1111111111111111111111111111111111111111111111111111111001011111;
MM[417] = 64'b1111111111111111111111111111111111111111111111111111111001011110;
MM[418] = 64'b1111111111111111111111111111111111111111111111111111111001011101;
MM[419] = 64'b1111111111111111111111111111111111111111111111111111111001011100;
MM[420] = 64'b1111111111111111111111111111111111111111111111111111111001011011;
MM[421] = 64'b1111111111111111111111111111111111111111111111111111111001011010;
MM[422] = 64'b1111111111111111111111111111111111111111111111111111111001011001;
MM[423] = 64'b1111111111111111111111111111111111111111111111111111111001011000;
MM[424] = 64'b1111111111111111111111111111111111111111111111111111111001010111;
MM[425] = 64'b1111111111111111111111111111111111111111111111111111111001010110;
MM[426] = 64'b1111111111111111111111111111111111111111111111111111111001010101;
MM[427] = 64'b1111111111111111111111111111111111111111111111111111111001010100;
MM[428] = 64'b1111111111111111111111111111111111111111111111111111111001010011;
MM[429] = 64'b1111111111111111111111111111111111111111111111111111111001010010;
MM[430] = 64'b1111111111111111111111111111111111111111111111111111111001010001;
MM[431] = 64'b1111111111111111111111111111111111111111111111111111111001010000;
MM[432] = 64'b1111111111111111111111111111111111111111111111111111111001001111;
MM[433] = 64'b1111111111111111111111111111111111111111111111111111111001001110;
MM[434] = 64'b1111111111111111111111111111111111111111111111111111111001001101;
MM[435] = 64'b1111111111111111111111111111111111111111111111111111111001001100;
MM[436] = 64'b1111111111111111111111111111111111111111111111111111111001001011;
MM[437] = 64'b1111111111111111111111111111111111111111111111111111111001001010;
MM[438] = 64'b1111111111111111111111111111111111111111111111111111111001001001;
MM[439] = 64'b1111111111111111111111111111111111111111111111111111111001001000;
MM[440] = 64'b1111111111111111111111111111111111111111111111111111111001000111;
MM[441] = 64'b1111111111111111111111111111111111111111111111111111111001000110;
MM[442] = 64'b1111111111111111111111111111111111111111111111111111111001000101;
MM[443] = 64'b1111111111111111111111111111111111111111111111111111111001000100;
MM[444] = 64'b1111111111111111111111111111111111111111111111111111111001000011;
MM[445] = 64'b1111111111111111111111111111111111111111111111111111111001000010;
MM[446] = 64'b1111111111111111111111111111111111111111111111111111111001000001;
MM[447] = 64'b1111111111111111111111111111111111111111111111111111111001000000;
MM[448] = 64'b1111111111111111111111111111111111111111111111111111111000111111;
MM[449] = 64'b1111111111111111111111111111111111111111111111111111111000111110;
MM[450] = 64'b1111111111111111111111111111111111111111111111111111111000111101;
MM[451] = 64'b1111111111111111111111111111111111111111111111111111111000111100;
MM[452] = 64'b1111111111111111111111111111111111111111111111111111111000111011;
MM[453] = 64'b1111111111111111111111111111111111111111111111111111111000111010;
MM[454] = 64'b1111111111111111111111111111111111111111111111111111111000111001;
MM[455] = 64'b1111111111111111111111111111111111111111111111111111111000111000;
MM[456] = 64'b1111111111111111111111111111111111111111111111111111111000110111;
MM[457] = 64'b1111111111111111111111111111111111111111111111111111111000110110;
MM[458] = 64'b1111111111111111111111111111111111111111111111111111111000110101;
MM[459] = 64'b1111111111111111111111111111111111111111111111111111111000110100;
MM[460] = 64'b1111111111111111111111111111111111111111111111111111111000110011;
MM[461] = 64'b1111111111111111111111111111111111111111111111111111111000110010;
MM[462] = 64'b1111111111111111111111111111111111111111111111111111111000110001;
MM[463] = 64'b1111111111111111111111111111111111111111111111111111111000110000;
MM[464] = 64'b1111111111111111111111111111111111111111111111111111111000101111;
MM[465] = 64'b1111111111111111111111111111111111111111111111111111111000101110;
MM[466] = 64'b1111111111111111111111111111111111111111111111111111111000101101;
MM[467] = 64'b1111111111111111111111111111111111111111111111111111111000101100;
MM[468] = 64'b1111111111111111111111111111111111111111111111111111111000101011;
MM[469] = 64'b1111111111111111111111111111111111111111111111111111111000101010;
MM[470] = 64'b1111111111111111111111111111111111111111111111111111111000101001;
MM[471] = 64'b1111111111111111111111111111111111111111111111111111111000101000;
MM[472] = 64'b1111111111111111111111111111111111111111111111111111111000100111;
MM[473] = 64'b1111111111111111111111111111111111111111111111111111111000100110;
MM[474] = 64'b1111111111111111111111111111111111111111111111111111111000100101;
MM[475] = 64'b1111111111111111111111111111111111111111111111111111111000100100;
MM[476] = 64'b1111111111111111111111111111111111111111111111111111111000100011;
MM[477] = 64'b1111111111111111111111111111111111111111111111111111111000100010;
MM[478] = 64'b1111111111111111111111111111111111111111111111111111111000100001;
MM[479] = 64'b1111111111111111111111111111111111111111111111111111111000100000;
MM[480] = 64'b1111111111111111111111111111111111111111111111111111111000011111;
MM[481] = 64'b1111111111111111111111111111111111111111111111111111111000011110;
MM[482] = 64'b1111111111111111111111111111111111111111111111111111111000011101;
MM[483] = 64'b1111111111111111111111111111111111111111111111111111111000011100;
MM[484] = 64'b1111111111111111111111111111111111111111111111111111111000011011;
MM[485] = 64'b1111111111111111111111111111111111111111111111111111111000011010;
MM[486] = 64'b1111111111111111111111111111111111111111111111111111111000011001;
MM[487] = 64'b1111111111111111111111111111111111111111111111111111111000011000;
MM[488] = 64'b1111111111111111111111111111111111111111111111111111111000010111;
MM[489] = 64'b1111111111111111111111111111111111111111111111111111111000010110;
MM[490] = 64'b1111111111111111111111111111111111111111111111111111111000010101;
MM[491] = 64'b1111111111111111111111111111111111111111111111111111111000010100;
MM[492] = 64'b1111111111111111111111111111111111111111111111111111111000010011;
MM[493] = 64'b1111111111111111111111111111111111111111111111111111111000010010;
MM[494] = 64'b1111111111111111111111111111111111111111111111111111111000010001;
MM[495] = 64'b1111111111111111111111111111111111111111111111111111111000010000;
MM[496] = 64'b1111111111111111111111111111111111111111111111111111111000001111;
MM[497] = 64'b1111111111111111111111111111111111111111111111111111111000001110;
MM[498] = 64'b1111111111111111111111111111111111111111111111111111111000001101;
MM[499] = 64'b1111111111111111111111111111111111111111111111111111111000001100;
MM[500] = 64'b1111111111111111111111111111111111111111111111111111111000001011;
MM[501] = 64'b1111111111111111111111111111111111111111111111111111111000001010;
MM[502] = 64'b1111111111111111111111111111111111111111111111111111111000001001;
MM[503] = 64'b1111111111111111111111111111111111111111111111111111111000001000;
MM[504] = 64'b1111111111111111111111111111111111111111111111111111111000000111;
MM[505] = 64'b1111111111111111111111111111111111111111111111111111111000000110;
MM[506] = 64'b1111111111111111111111111111111111111111111111111111111000000101;
MM[507] = 64'b1111111111111111111111111111111111111111111111111111111000000100;
MM[508] = 64'b1111111111111111111111111111111111111111111111111111111000000011;
MM[509] = 64'b1111111111111111111111111111111111111111111111111111111000000010;
MM[510] = 64'b1111111111111111111111111111111111111111111111111111111000000001;
MM[511] = 64'b0111111111111111111111111111111111111111111111111111111000000000;
end
Select S(MM[t],bo,temp);

always @(x)
begin
	
	if(tag[0] == t)
	begin
		flag <= 1;
		index <= 0;
	end

	if(tag[1] == t)
	begin
		flag <= 1;
		index <= 1;	
	end

	if(tag[2] == t)
	begin
		flag <= 1;
		index <= 2;	
	end

	if(tag[3] == t)
	begin
		flag <= 1;
		index <= 3;	
	end

	if(tag[4] == t)
	begin
		flag <= 1;
		index <= 4;	
	end

	if(tag[5] == t)
	begin
		flag <= 1;
		index <= 5;	
	end

	if(tag[6] == t)
	begin
		flag <= 1;
		index <= 6;	
	end	

	if(tag[7] == t)
	begin
		flag <= 1;
		index <= 7;	
	end

	if(flag == 1)
	begin	
		y <= 1'b1;
	end

	else
		begin	
			y <= 1'b0;
			cache[pointer] <= MM[t];
			tag[pointer] <= t;
			pointer = pointer + 1;
		end
end
assign word = temp;
assign counter = pointer;
endmodule